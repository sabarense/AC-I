module exercicio_04(input [7:0] num_bin, output [7:0] resultado);
  assign resultado = num_bin * 4; // Parte b)
endmodule
